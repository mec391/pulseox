module frame_storage( 
//this module receives data from the the ALU, 
//determines what the frame should be, 
//and sends frames to the the TFT driver pixel by pixel


);


endmodule